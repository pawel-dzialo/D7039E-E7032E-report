** Profile: "SCHEMATIC1-sweep"  [ C:\Cadence\Projects\Skola\Projektkurs\Antialiasing-PSpiceFiles\SCHEMATIC1\sweep.sim ] 

** Creating circuit file "sweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "C:\Cadence\Projects\Projekt174\Libary\ad711.lib" 
.lib "C:\Cadence\SPB_17.4\tools\pspice\library\opamp.lib" 
.lib "C:\Cadence\LTU_Parts\LTU10.LIB" 
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 1 10k
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
