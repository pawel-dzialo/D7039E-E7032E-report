** Profile: "IdealOPamp-transientGain"  [ c:\cadence\projects\skola\projektkurs\eeg_amplifier-pspicefiles\idealopamp\transientgain.sim ] 

** Creating circuit file "transientGain.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../eeg_amplifier-pspicefiles/opamp_int.lib" 
.LIB "../../../eeg_amplifier-pspicefiles/eeg_amplifier.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "C:\Cadence\Projects\Projekt174\Libary\ad711.lib" 
.lib "C:\Cadence\SPB_17.4\tools\pspice\library\opamp.lib" 
.lib "C:\Cadence\LTU_Parts\LTU10.LIB" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 0.05 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\IdealOPamp.net" 


.END
